`timescale 1ns / 1ns

// verilator lint_off UNUSED
// verilator lint_off UNDRIVEN

module blk_mem_gen_1
    (
        input wire [8:0] addra,
        input wire clka,
        output wire [63:0] douta
    );
endmodule

// verilator lint_on UNUSED
// verilator lint_on UNDRIVEN
