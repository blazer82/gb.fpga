`timescale 1ns / 1ns

// verilator lint_off UNUSED
// verilator lint_off UNDRIVEN

module clk_wiz_0
    (
        input wire clk_in1,
        output wire clk_out1,
        output wire clk_out2
    );
endmodule

// verilator lint_on UNUSED
// verilator lint_on UNDRIVEN
