`timescale 1ns / 1ns

module STARTUPE2
    #(
        parameter PROG_USR = "FALSE",
        parameter SIM_CCLK_FREQ = 0.0
    )
    (
        input wire GSR,
        input wire GTS,
        input wire USRCCLKO,
        input wire USRCCLKTS,
        input wire USRDONEO
    );
endmodule
