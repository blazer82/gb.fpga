`timescale 1ns / 1ns

module clk_wiz_0
    (
        input wire clk_in1,
        output wire clk_out1,
        output wire clk_out2
    );
endmodule
