`timescale 1ns / 1ns

module blk_mem_gen_1
    (
        input wire [8:0] addra,
        input wire clka,
        output wire [63:0] douta
    );
endmodule
